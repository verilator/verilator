// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2020 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

class Cls1;
   function int randomize;
      return 1;
   endfunction
endclass

class Cls2;
   function void randomize(int x);
   endfunction
   function void srandom(int seed);
   endfunction
endclass

module t;
endmodule
