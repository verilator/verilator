// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2024 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

// Rather than look at waivers, just check we included it
`ifndef _VERILATED_STD_WAIVER_VLT_
`error "Didn't include, no _VERILATED_STD_WAIVER_VLT_"
`endif

module t;
endmodule
