module top (
   input logic[26:72][52:73][123:33][3:42] multidim_signal
);
endmodule
