// DESCRIPTION: Verilator: Large test for SystemVerilog

// This file ONLY is placed under the Creative Commons Public Domain, for
// SPDX-FileCopyrightText: 2012
// SPDX-License-Identifier: CC0-1.0

// Contributed by M W Lund, Atmel Corporation.

//*****************************************************************************
// PAD_GND - Ground Supply Pad (Dummy!!!!)
//*****************************************************************************

module pad_gnd
#( parameter ID = 0 )
  (
   inout wire pad
   );

  assign pad = 1'b0;
endmodule // pad_gnd
