// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2023 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

class Packet;
   rand int one;

   constraint a { one > 0 && one < 2; }

   constraint empty { }

endclass

module t;

   Packet p;

   int v;

   initial begin
      p = new;
      v = p.randomize();
      if (v != 1) $stop;
      if (p.one != 1) $stop;

      $write("*-* All Finished *-*\n");
      $finish;
   end
endmodule
