// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2022 by Antmicro Ltd.
// SPDX-License-Identifier: CC0-1.0

module t (/*AUTOARG*/);
   reg [3:0] a = 4'b11z1;
   logic     b = 1'z === a[1];
   always begin
      if (b) begin
         $write("*-* All Finished *-*\n");
         $finish;
      end
   end
endmodule
