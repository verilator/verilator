// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2009 by Wilson Snyder.

module t;
   reg foobar;

   task boobar; endtask

   initial begin
      if (foobat) $stop;
      boobat;
   end
endmodule
