// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2025 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;

   typedef int arr_t [5];
   arr_t arr;
   localparam type arr_type = type(arr);
   arr_type arr_prime;

   initial begin
      arr[3] = 123;
      arr_prime = arr;
      if (arr_prime[3] != 123) $stop();
      $write("*-* All Finished *-*\n");
      $finish;
   end

endmodule
