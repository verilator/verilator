// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2019 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;
   initial begin
      int i;

      i = {} + 1;

      i = {};

      $write("*-* All Finished *-*\n");
      $finish;
   end
endmodule
