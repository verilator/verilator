
interface bus_if #(
   parameter int p_awidth = 4
   ,parameter int p_dwidth = 7
);
   typedef struct packed {
      logic [p_awidth-1:0] addr;
   } rq_t;
   typedef struct packed {
      logic [p_dwidth-1:0] data;
   } rs_t;

   rq_t rq;
   rs_t rs;
endinterface

module a_mod(
   bus_if bus_io
);
   localparam bus_rq_t = bus_io.rq_t;
   localparam bus_rs_t = bus_io.rs_t;
   localparam p_awidth = bus_io.p_awidth;
   localparam p_dwidth = bus_io.p_dwidth;

   bus_rq_t rq;
   bus_rs_t rs;

   assign rs.data = 8'ha5;
   assign bus_io.rs = rs;

endmodule

module top();
   bus_if #(.p_awidth(16), .p_dwidth(8)) bus_io();

   a_mod a_mod_inst(
      .bus_io(bus_io)
   );

   initial begin
      #1;
      if(bus_io.rs.data != 8'ha5) $stop;
      $write("*-* All Finished *-*\n");
      $finish;
   end
endmodule
