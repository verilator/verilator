// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2019 by Wilson Snyder.

module t (/*AUTOARG*/);

   int u1;
   int u1;
   int u1;
   int u1;
   int u1;
   int u1;
   int u1;

endmodule
