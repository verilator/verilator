// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2024 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

class Cls#(type T = bit);
endclass

module t;

   Cls#(bit) cb;

   Cls#(Cls#(bit)) ccb;

   initial begin
      $write("*-* All Finished *-*\n");
      $finish;
   end

endmodule
