// DESCRIPTION: Verilator: Verilog dummy test module
//
// This file ONLY is placed under the Creative Commons Public Domain
// SPDX-FileCopyrightText: 2022 Yu-Sheng Lin
// SPDX-License-Identifier: CC0-1.0

module t(input clk);
endmodule
