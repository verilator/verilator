// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2014 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;

   string s;
   integer i;

   // Check constification
   initial begin
      s="1234";
      i = s.len(0); // BAD
      s.itoa;  // BAD
      s.itoa(1,2,3);  // BAD
      s.bad_no_such_method();  // BAD
   end

endmodule
