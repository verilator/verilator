// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2023 Antmicro Ltd
// SPDX-License-Identifier: CC0-1.0

module t;
   initial begin
      int q[5];

      q.mex;

      $write("*-* All Finished *-*\n");
      $finish;
   end
endmodule
