// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2014 by Wilson Snyder.

`define checkh(gotv,expv) do if ((gotv) !== (expv)) begin $write("%%Error: %s:%0d:  got='h%x exp='h%x\n", `__FILE__,`__LINE__, (gotv), (expv)); $stop; end while(0);
`define checks(gotv,expv) do if ((gotv) !== (expv)) begin $write("%%Error: %s:%0d:  got='%s' exp='%s'\n", `__FILE__,`__LINE__, (gotv), (expv)); $stop; end while(0);

module t (/*AUTOARG*/
   // Inputs
   clk
   );
   input clk;

   logic [2:0] foo [1:0];
   initial begin
      foo[0] = 3'b101;
      foo[1] = 3'b011;

      `checkh(foo.or, 3'b111);
      `checkh(foo.and, 3'b001);
      `checkh(foo.xor, 3'b110);

      $write("*-* All Finished *-*\n");
      $finish;
   end

endmodule
