// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2022 Antmicro Ltd
// SPDX-License-Identifier: CC0-1.0

module t(/*AUTOARG*/
   // Inputs
   rstn
   );
   input rstn;

   default disable iff (!rstn);
   default disable iff (!rstn);

endmodule
