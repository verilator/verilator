// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2009 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

module t;
   reg foobar;

   task boobar; endtask

   initial begin
      if (foobat) $stop;
      boobat;
   end
endmodule
