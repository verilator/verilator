// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2003 by Wilson Snyder.

typedef enum { HIDE_VALUE = 0 } hide_enum_t;

module t;

   typedef enum { HIDE_VALUE = 0 } hide_enum_t;

endmodule
