// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2025 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

// 6.21 Scope and lifetime
// Automatic variables and elements of dynamically sized array variables shall
// not be written with nonblocking, continuous, or procedural continuous
// assignments. Non-static class properties shall not be written with continuous
// or procedural continuous assignments.

class Cls;
  static int s_ok1;
  static int s_ok2;
  int m_bad1;
  int m_bad2;
endclass

module t(clk);
  input clk;

  Cls c;

  automatic int bad_auto3;
  automatic int bad_auto4;
  int bad_dyn5[];
  int bad_dyn6[];
  int empty_dyn[];

  assign bad_auto3 = 2;  // <--- Error: continuous automatic
  assign bad_dyn5 = empty_dyn;  // <--- Error: continuous dynarray
  assign c.m_bad1 = 2;  // <--- Error: continuous class non-static
  // Only one simulator fails on this, probably not legal
  // assign Cls::s_ok1 = 2;  // OK: continuous class static

  logic ok_7;
  task mt(output o);  // OK: function output
    o <= 1;
  endtask

  always @(posedge clk) begin
    bad_auto4 <= 2;  // <--- Error: nonblocking automatic
    bad_dyn6 <= empty_dyn;  // <--- Error: nonblocking dynarray
    Cls::s_ok2 <= 2;  // OK: nonblocking class static
    c.m_bad2 <= 2;  // <--- Error: nonblocking class automatic
    mt(ok_7);
    $stop;
  end

endmodule
