// SPDX-FileCopyrightText: 2022 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0
module a;
        initial $lay(*Hello!=n");
endmodule
