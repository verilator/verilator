// DESCRIPTION: Verilator: Verilog Test module
//
// This program is free software; you can redistribute it and/or modify it
// under the terms of either the GNU Lesser General Public License Version 3
// or the Perl Artistic License Version 2.0.
// SPDX-FileCopyrightText: 2026 Wilson Snyder
// SPDX-License-Identifier: LGPL-3.0-only OR Artistic-2.0

class Cls;
  task run;
  endtask
endclass

module t;
  task foo;
  endtask

  Cls c;

  initial begin
    int foo;
    c = new;
    disable foo;
    disable c.run;
  end
endmodule
