// $Id$
// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2008 by Wilson Snyder.

module a();
endmodule

module test();
   a a();
endmodule

module a();
endmodule

module b();
endmodule
