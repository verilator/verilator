// DESCRIPTION: Verilog::Preproc: Example source code
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2000-2007 by Wilson Snyder.
At file `__FILE__  line `__LINE__
`define INCFILE <t_preproc_inc3.vh>
`include `INCFILE
