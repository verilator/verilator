// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2010 by Wilson Snyder.

//See bug289

`include "t_preproc_inc_inc_bad.vh"

module t;
endmodule
