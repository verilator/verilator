// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2012 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

module t;
   initial Pkg::hello();  //<--- Warning
endmodule
package Pkg;
   function void hello(); endfunction
endpackage
