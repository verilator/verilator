// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2003 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

typedef enum { HIDE_VALUE = 0 } hide_enum_t;

module t;

   typedef enum { HIDE_VALUE = 0 } hide_enum_t;

endmodule
