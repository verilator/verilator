// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2026 by Antmicro.
// SPDX-License-Identifier: CC0-1.0

module t;
  sub \x.y  ();
  initial begin
    $write("*-* All finished *-*\n");
    $finish;
  end
endmodule

module sub;
        bit z;
endmodule

