// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2019 by Wilson Snyder.

// Legal with ANSI Verilog 2001 style ports
module t
  (
   output wire ok_ow,
   output reg  ok_or);

   wire ok_o_w;
   reg   ok_o_r;
endmodule
