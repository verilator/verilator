// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2019 by Wilson Snyder.

module t (/*AUTOARG*/);

<<<<<<< HEAD  // Intentional test: This conflict marker should be here
   initial $display("Hello");
=======   // Intentional test: This conflict marker should be here
   initial $display("Goodbye");
>>>>>>> MERGE  // Intentional test: This conflict marker should be here

endmodule
