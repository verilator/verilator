// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2010 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

inc line 6;
inc line 7;  // example_lint_off_line FOO
inc line 8;  // example_lint_off_line BAR
inc line 9;
