// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2020 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

module t;

   integer a[];

   string  s;

   initial begin
      s = "str";
      a = new [s];  // Bad
   end

endmodule
