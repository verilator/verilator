module t();
    reg x;
/* verilator public_off */
endmodule
