// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2024 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

class Packet;
   extern constraint missing_bad;
endclass

constraint Packet::missing_extern { }

module t (/*AUTOARG*/);
endmodule
