// ======================================================================
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty.
// SPDX-License-Identifier: CC0-1.0
// ======================================================================

module t;
  logic unpacked[1]  /*verilator forceable*/;
endmodule
