// DESCRIPTION: Verilog::Preproc: Example source code
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2000-2007 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0
At file `__FILE__  line `__LINE__
`define INCFILE <t_preproc_inc3.vh>
`include `INCFILE
