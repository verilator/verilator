// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2003 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;
   string s = "a string";
   initial begin
      $display("%d %x %f %t", s, s, s, s);
      $write("*-* All Finished *-*\n");
      $finish;
   end
endmodule
