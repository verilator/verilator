// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2019 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;

<<<<<<< HEAD  // Intentional test: This conflict marker should be here
   initial $display("Hello");
=======   // Intentional test: This conflict marker should be here
   initial $display("Goodbye");
>>>>>>> MERGE  // Intentional test: This conflict marker should be here

endmodule
