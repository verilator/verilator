// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2016 by Wilson Snyder.

module t
   (
   input wire rst
   );

   integer q;
   
   always @(*)
     if (rst)
       assign q = 0;
     else
       deassign q;

endmodule
