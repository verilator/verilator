// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2023 Anthony Donlon
// SPDX-License-Identifier: CC0-1.0

module t;
    m ();
    m ();
endmodule

module m;
endmodule
