// DESCRIPTION: Verilator: Verilog dummy test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2022 by Yu-Sheng Lin.
// SPDX-License-Identifier: CC0-1.0

module t(input clk);
endmodule
