// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2018 by Wilson Snyder.

package defs;
   int sig;
endpackage

import defs::*;

module t;
endmodule
