// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2025 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

`include "t_flag_f_tsub_inc.v"

`ifndef GOT_DEF5
`error "No GOT_DEF5"
`endif

module t;
endmodule
