// DESCRIPTION: Verilator: Verilog Test module

module t;
   initial begin
      // verilator lint_off FUTURE1
      $write("*-* All Finished *-*\n");
      $finish;
      // verilator FUTURE2
      // verilator FUTURE2 blah blah
   end
endmodule
