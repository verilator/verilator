// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2020 by Wilsn Snyder.
// SPDX-License-Identifier: CC0-1.0

module t
  (
   output id0
   );

   assign id0 = 0;

endmodule
