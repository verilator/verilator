// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2011 by Wilson Snyder.

module sub;
   integer i;
   initial begin
      i = 23.2;
   end
endmodule
