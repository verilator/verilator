module a;
	initial $lay(*Hello!=n");
endmodule
