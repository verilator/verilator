// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2005-2007 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;

   parameter [200:0] MIXED = 32'dx_1;

endmodule
