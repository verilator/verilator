// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2025 by Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

package pkg;
endpackage

class genericClass;
  import pkg::*;
endclass

module tb_top ();
endmodule
