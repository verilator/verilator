// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2024 by Antmicro.
// SPDX-License-Identifier: CC0-1.0

`define DISPLAY_PASS(file, line) \
   $display("Passed '%m' at %s:%g", file, line)

`define DISPLAY_FAIL(file, line) \
   $display("Failed '%m' at %s:%g", file, line)

`define RUN_ALL_ASSERTS \
   $display("==========\nRunning all asserts at: %s:%g\n==========", `__FILE__, `__LINE__); \
   run_all_asserts(`__FILE__, `__LINE__); \
   cover_simple_immediate_`__LINE__: cover(0); \
   cover_simple_immediate_stmt_`__LINE__: cover(0) `DISPLAY_PASS(`__FILE__, `__LINE__); \
   cover_observed_deferred_immediate_`__LINE__: cover #0 (0); \
   cover_observed_deferred_immediate_stmt_`__LINE__: cover #0 (0) `DISPLAY_PASS(`__FILE__, `__LINE__); \
   cover_final_deferred_immediate_`__LINE__: cover final (0); \
   cover_final_deferred_immediate_stmt_`__LINE__: cover final (0) `DISPLAY_PASS(`__FILE__, `__LINE__); \

module t (/*AUTOARG*/
   clk
   );
   input clk;

   let ON = 3;
   let OFF = 4;
   let KILL = 5;

   let CONCURRENT = 1; 
   let SIMPLE_IMMEDIATE = 2;
   let OBSERVED_DEFERRED_IMMEDIATE = 4;
   let FINAL_DEFERRED_IMMEDIATE = 8;
   let UNIQUE = 32;
   let UNIQUE0 = 64;
   let PRIORITY = 128;

   let ALL = 255;

   /* CONCURRENT|SIMPLE_IMMEDIATE|OBSERVED_DEFERRED_IMMEDIATE|FINAL_DEFERRED_IMMEDIATE */
   let ALL_ASSERTIONS = 15;

   concurrent concurrent(.clk(clk));

   initial begin
      // simple immediate
      $assertcontrol(OFF, ALL);
      $assertcontrol(ON, SIMPLE_IMMEDIATE);
      `RUN_ALL_ASSERTS
      $assertcontrol(OFF, SIMPLE_IMMEDIATE);
      `RUN_ALL_ASSERTS

      // observed deferred immediate
      $assertcontrol(OFF, ALL);
      $assertcontrol(ON, OBSERVED_DEFERRED_IMMEDIATE);
      `RUN_ALL_ASSERTS
      $assertcontrol(OFF, OBSERVED_DEFERRED_IMMEDIATE);
      `RUN_ALL_ASSERTS

      // final deferred immediate
      $assertcontrol(OFF, ALL);
      $assertcontrol(ON, FINAL_DEFERRED_IMMEDIATE);
      `RUN_ALL_ASSERTS
      $assertcontrol(OFF, FINAL_DEFERRED_IMMEDIATE);
      `RUN_ALL_ASSERTS

      // on, off, kill test
      $assertoff;
      `RUN_ALL_ASSERTS;
      $asserton;
      `RUN_ALL_ASSERTS;
      $assertkill;
      `RUN_ALL_ASSERTS;

      $assertcontrol(ON, 6 /*SIMPLE_IMMEDIATE | OBSERVED_DEFERRED_IMMEDIATE*/);
      `RUN_ALL_ASSERTS;
      $assertcontrol(ON, FINAL_DEFERRED_IMMEDIATE);
      `RUN_ALL_ASSERTS;
      $assertcontrol(OFF, 12 /*OBSERVED_DEFERRED_IMMEDIATE|FINAL_DEFERRED_IMMEDIATE*/);
      `RUN_ALL_ASSERTS;
      $assertcontrol(OFF, FINAL_DEFERRED_IMMEDIATE);
      `RUN_ALL_ASSERTS;
      $assertcontrol(OFF, SIMPLE_IMMEDIATE);
      `RUN_ALL_ASSERTS;
      $assertcontrol(ON, SIMPLE_IMMEDIATE);
      `RUN_ALL_ASSERTS;
      $assertcontrol(OFF, ALL);
      `RUN_ALL_ASSERTS;
      $assertcontrol(ON, ALL);
      `RUN_ALL_ASSERTS;
      $assertcontrol(KILL, ALL);
      `RUN_ALL_ASSERTS;
      $assertcontrol(ON, ALL_ASSERTIONS);
      `RUN_ALL_ASSERTS;
      $assertcontrol(OFF, ALL_ASSERTIONS);
      `RUN_ALL_ASSERTS;

      // concurrent test
      #10;
      $display("Disabling concurrent asserts, time: %g", $time);
      $assertcontrol(ON, ALL);
      $assertcontrol(OFF, CONCURRENT);
      #10;
      $display("Enabling concurrent asserts, time: %g", $time);
      $assertcontrol(ON, CONCURRENT);
      $finish;
   end
endmodule

task run_all_asserts(string file, integer line);
   run_simple_immediate(file, line);
   run_observed_deferred_immediate(file, line);
   run_final_deferred_immediate(file, line);
   // TODO
   //run_if_case(file, line);
endtask

task run_simple_immediate(string file, integer line);
   $display("Testing assert_simple_immediate at %s:%g", file, line);
   assert_simple_immediate: assert(0);
   assert_simple_immediate_else: assert(0) else `DISPLAY_FAIL(file, line);
   assert_simple_immediate_stmt: assert(0) `DISPLAY_PASS(file, line);
   assert_simple_immediate_stmt_else: assert(0) `DISPLAY_PASS(file, line); else `DISPLAY_FAIL(file, line);

   $display("Testing assume_simple_immediate at %s:%g", file, line);
   assume_simple_immediate: assume(0);
   assume_simple_immediate_else: assume(0) else `DISPLAY_FAIL(file, line);
   assume_simple_immediate_stmt: assume(0) `DISPLAY_PASS(file, line);
   assume_simple_immediate_stmt_else: assume(0) `DISPLAY_PASS(file, line); else `DISPLAY_FAIL(file, line);
endtask

task run_observed_deferred_immediate(string file, integer line);
   $display("Testing assert_observed_deferred_immediate at %s:%g", file, line);
   assert_observed_deferred_immediate: assert #0 (0);
   assert_observed_deferred_immediate_else: assert #0 (0) else `DISPLAY_FAIL(file, line);
   assert_observed_deferred_immediate_stmt: assert #0 (0) `DISPLAY_PASS(file, line);
   assert_observed_deferred_immediate_stmt_else: assert #0 (0) `DISPLAY_PASS(file, line); else `DISPLAY_FAIL(file, line);

   $display("Testing assume_observed_deferred_immediate at %s:%g", file, line);
   assume_observed_deferred_immediate: assume #0 (0);
   assume_observed_deferred_immediate_else: assume #0 (0) else `DISPLAY_FAIL(file, line);
   assume_observed_deferred_immediate_stmt: assume #0 (0) `DISPLAY_PASS(file, line);
   assume_observed_deferred_immediate_stmt_else: assume #0 (0) `DISPLAY_PASS(file, line); else `DISPLAY_FAIL(file, line);
endtask

task run_final_deferred_immediate(string file, integer line);
   $display("Testing assert_final_deferred_immediate at %s:%g", file, line);
   assert_final_deferred_immediate: assert final (0);
   assert_final_deferred_immediate_else: assert final (0) else `DISPLAY_FAIL(file, line);
   assert_final_deferred_immediate_stmt: assert final (0) `DISPLAY_PASS(file, line);
   assert_final_deferred_immediate_stmt_else: assert final (0) `DISPLAY_PASS(file, line); else `DISPLAY_FAIL(file, line);

   $display("Testing assume_final_deferred_immediate at %s:%g", file, line);
   assume_final_deferred_immediate: assume final (0);
   assume_final_deferred_immediate_else: assume final (0) else `DISPLAY_FAIL(file, line);
   assume_final_deferred_immediate_stmt: assume final (0) `DISPLAY_PASS(file, line);
   assume_final_deferred_immediate_stmt_else: assume final (0) `DISPLAY_PASS(file, line); else `DISPLAY_FAIL(file, line);
endtask

task run_if_case(string file, integer line);
   $display("Testing unique0_if at %s:%g", file, line);
   unique0_if: unique0 if (0) `DISPLAY_PASS(file, line);
   unique0_if_else: unique0 if (0) `DISPLAY_PASS(file, line); else `DISPLAY_FAIL(file, line);
   $display("Testing unique_if at %s:%g", file, line);
   unique_if: unique if (0) `DISPLAY_PASS(file, line);
   unique_if_else: unique if (0) `DISPLAY_PASS(file, line); else `DISPLAY_FAIL(file, line);
   $display("Testing priority_if at %s:%g", file, line);
   priority_if: priority if (0) `DISPLAY_PASS(file, line);
   priority_if_else: priority if (0) `DISPLAY_PASS(file, line); else `DISPLAY_FAIL(file, line);

   $display("Testing unique0_case at %s:%g", file, line);
   unique0_case: unique0 case (0) 1: `DISPLAY_PASS(file, line); endcase
   unique0_case_default: unique0 case (0) 1: `DISPLAY_PASS(file, line); default: `DISPLAY_FAIL(file, line); endcase
   $display("Testing unique_case at %s:%g", file, line);
   unique_case: unique case (0) 1: `DISPLAY_PASS(file, line); endcase
   unique_case_default: unique case (0) 1: `DISPLAY_PASS(file, line); default: `DISPLAY_FAIL(file, line); endcase
   $display("Testing priority_case at %s:%g", file, line);
   priority_case: priority case (0) 1: `DISPLAY_PASS(file, line); endcase
   priority_case_default: priority case (0) 1: `DISPLAY_PASS(file, line); default: `DISPLAY_FAIL(file, line); endcase
endtask

module concurrent(input clk);
   property prop();
      @(posedge clk) 0
   endproperty

   assert_concurrent: assert property (prop);
   assert_concurrent_else: assert property(prop) else `DISPLAY_FAIL(`__FILE__, `__LINE__);
   assert_concurrent_stmt: assert property(prop) `DISPLAY_PASS(`__FILE__, `__LINE__);
   assert_concurrent_stmt_else: assert property(prop) `DISPLAY_PASS(`__FILE__, `__LINE__); else `DISPLAY_FAIL(`__FILE__, `__LINE__);

   assume_concurrent: assume property(prop);
   assume_concurrent_else: assume property(prop) else `DISPLAY_FAIL(`__FILE__, `__LINE__);
   assume_concurrent_stmt: assume property(prop) `DISPLAY_PASS(`__FILE__, `__LINE__);
   assume_concurrent_stmt_else: assume property(prop) `DISPLAY_PASS(`__FILE__, `__LINE__); else `DISPLAY_FAIL(`__FILE__, `__LINE__);

   cover_concurrent: cover property(prop);
   cover_concurrent_stmt: cover property(prop) `DISPLAY_PASS(`__FILE__, `__LINE__);
endmodule
