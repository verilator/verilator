// DESCRIPTION: Verilator: Verilog Test module
//
// Copyright 2020 by Wilson Snyder. This program is free software; you can
// redistribute it and/or modify it under the terms of either the GNU
// Lesser General Public License Version 3 or the Perl Artistic License
// Version 2.0.

module t;
   export "DPI-C" task dpix_task;
   task dpix_task();
      $write("Hello in %m\n");
   endtask
endmodule
