// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2020 by Dan Petrisko.
// SPDX-License-Identifier: CC0-1.0

typedef struct packed {
   logic clk /*verilator clocker*/;
   logic data;
} ss_s;

endmodule
