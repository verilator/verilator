module t;

endmodule
