// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2017 by Wilson Snyder.

module t (input mispkg::foo_t a);
   reg mispkgb::bar_t b;
endmodule
