// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2005 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;

   looped looped ();

endmodule

module looped;
   looped2 looped2 ();
endmodule

module looped2;
   looped looped ();
endmodule
