// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2019 by Wilson Snyder.

module t_multitop1s;
   initial $display("In '%m'");
endmodule

module in_subfile;
   initial $display("In '%m'");
endmodule
