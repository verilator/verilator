module t_emit_accessors(
    input bit a,
    output bit b
);

endmodule;