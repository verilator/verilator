// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2020 by Edgar E. Iglesias.
// SPDX-License-Identifier: CC0-1.0

module t (
   clk
   );
   input clk;
endmodule
