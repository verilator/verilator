// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2017 by Wilson Snyder.

module t;
   bit [256:0] num = 'd123456789123456789123456789;
endmodule
