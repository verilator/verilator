// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2022 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;

   int array[2][2];

   initial begin
      foreach (array[i, j, badk, badl]);  // bad

      $stop;
   end

endmodule
