// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2024 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

// Rather than look at waivers, just check we included it
`ifdef _VERILATED_STD_WAIVER_VLT_
`error "Shouldn't have included _VERILATED_STD_WAIVER_VLT_"
`endif

module t;
endmodule
