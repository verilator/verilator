// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2020 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

/* verilator lint_off PINNOTFOUND */
module a;
localparam A=1;
generate
if (A==0)
begin
b b_inst(.x(1'b0));
end
endgenerate
endmodule

module b;
endmodule
