// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2024 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

module t(/*AUTOARG*/);
   defparam id_13.id_14 = -id_13,
     id_15 = id_14;

   defparam id_8 = 1, id_9 = 1;
endmodule
