// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2023 Antmicro Ltd
// SPDX-License-Identifier: CC0-1.0

class Foo#(type T = logic) extends T;
endclass

module t;
   initial begin
      $write("*-* All Finished *-*\n");
      $finish;
   end
endmodule
