// $Id:$
// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2003 by Wilson Snyder.

module t (/*AUTOARG*/
   // Inputs
   clk
   );
   parameter PAR = 3;
   input clk;

   defparam i.L00 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L01 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L02 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L03 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L04 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L05 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L06 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L07 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L08 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L09 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L0A = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L0B = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L0C = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L0D = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L0E = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L0F = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L10 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L11 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L12 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L13 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L14 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L15 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L16 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L17 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L18 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L19 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L1A = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L1B = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L1C = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L1D = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L1E = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L1F = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L20 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L21 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L22 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L23 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L24 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L25 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L26 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L27 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L28 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L29 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L2A = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L2B = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L2C = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L2D = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L2E = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L2F = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L30 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L31 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L32 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L33 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L34 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L35 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L36 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L37 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L38 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L39 = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L3A = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L3B = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L3C = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L3D = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L3E = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.L3F = 256'h000012300000000000000000000000000000000000000000000000000000cdef;
   defparam i.A0 = "HELLO_WORLD_BOY_THIS_IS_LONG";
   defparam i.A1 = "HELLO_WORLD_BOY_THIS_IS_LONG";
   defparam i.A2 = "HELLO_WORLD_BOY_THIS_IS_LONG";

   i i (.clk(clk));

   integer cyc=1;
   always @ (posedge clk) begin
      cyc <= cyc + 1;
      if (cyc==1) begin
	 $write("*-* All Finished *-*\n");
	 $finish;
      end
   end

endmodule

module i
    (/*AUTOARG*/
   // Inputs
   clk
   );

   // verilator public_module

   input       clk;

   parameter [255:0] L00 = 256'h0;
   parameter [255:0] L01 = 256'h0;
   parameter [255:0] L02 = 256'h0;
   parameter [255:0] L03 = 256'h0;
   parameter [255:0] L04 = 256'h0;
   parameter [255:0] L05 = 256'h0;
   parameter [255:0] L06 = 256'h0;
   parameter [255:0] L07 = 256'h0;
   parameter [255:0] L08 = 256'h0;
   parameter [255:0] L09 = 256'h0;
   parameter [255:0] L0A = 256'h0;
   parameter [255:0] L0B = 256'h0;
   parameter [255:0] L0C = 256'h0;
   parameter [255:0] L0D = 256'h0;
   parameter [255:0] L0E = 256'h0;
   parameter [255:0] L0F = 256'h0;
   parameter [255:0] L10 = 256'h0;
   parameter [255:0] L11 = 256'h0;
   parameter [255:0] L12 = 256'h0;
   parameter [255:0] L13 = 256'h0;
   parameter [255:0] L14 = 256'h0;
   parameter [255:0] L15 = 256'h0;
   parameter [255:0] L16 = 256'h0;
   parameter [255:0] L17 = 256'h0;
   parameter [255:0] L18 = 256'h0;
   parameter [255:0] L19 = 256'h0;
   parameter [255:0] L1A = 256'h0;
   parameter [255:0] L1B = 256'h0;
   parameter [255:0] L1C = 256'h0;
   parameter [255:0] L1D = 256'h0;
   parameter [255:0] L1E = 256'h0;
   parameter [255:0] L1F = 256'h0;
   parameter [255:0] L20 = 256'h0;
   parameter [255:0] L21 = 256'h0;
   parameter [255:0] L22 = 256'h0;
   parameter [255:0] L23 = 256'h0;
   parameter [255:0] L24 = 256'h0;
   parameter [255:0] L25 = 256'h0;
   parameter [255:0] L26 = 256'h0;
   parameter [255:0] L27 = 256'h0;
   parameter [255:0] L28 = 256'h0;
   parameter [255:0] L29 = 256'h0;
   parameter [255:0] L2A = 256'h0;
   parameter [255:0] L2B = 256'h0;
   parameter [255:0] L2C = 256'h0;
   parameter [255:0] L2D = 256'h0;
   parameter [255:0] L2E = 256'h0;
   parameter [255:0] L2F = 256'h0;
   parameter [255:0] L30 = 256'h0;
   parameter [255:0] L31 = 256'h0;
   parameter [255:0] L32 = 256'h0;
   parameter [255:0] L33 = 256'h0;
   parameter [255:0] L34 = 256'h0;
   parameter [255:0] L35 = 256'h0;
   parameter [255:0] L36 = 256'h0;
   parameter [255:0] L37 = 256'h0;
   parameter [255:0] L38 = 256'h0;
   parameter [255:0] L39 = 256'h0;
   parameter [255:0] L3A = 256'h0;
   parameter [255:0] L3B = 256'h0;
   parameter [255:0] L3C = 256'h0;
   parameter [255:0] L3D = 256'h0;
   parameter [255:0] L3E = 256'h0;
   parameter [255:0] L3F = 256'h0;
   parameter [255:0] A0 = 256'h0;
   parameter [255:0] A1 = 256'h0;
   parameter [255:0] A2 = 256'h0;

   always @ (posedge clk) begin
   end
endmodule
