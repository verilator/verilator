// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2010 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

module t
   (
  input wire i,
  input wire i2 = i   // Good under IEEE 1800-2009
   );

endmodule
