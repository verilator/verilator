// DESCRIPTION: Verilator: Verilog example module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2017 by Wilson Snyder.

// See also the EXAMPLE section in the verilator manpage/document.
module top;
   initial begin
      $display("Hello World!");
      $finish;
   end
endmodule
