/* verilator public_on */
/* verilator public_on */
module t();
    reg x;
endmodule
/* verilator public_off */