// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2020 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0
//

module t (/*AUTOARG*/);

   class Cls;

      static task static_task();
      endtask

   endclass : Cls

   initial begin
      Cls::static_task();
      $finish;
   end

endmodule
