// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2007 by Wilson Snyder.

module t (/*AUTOARG*/
   // Outputs
   ok, o, og, org,
   // Inputs
   i
   );

   reg    a;
   reg    a;

   integer l;
   integer l;

   bit     b;
   bit     b;

   output ok;
   reg    ok;

   output o;
   output o;

   input  i;
   input  i;

   output oi;
   input  oi;

   output og;
   reg    og;
   reg    og;

   output reg org;
   output reg org;

endmodule
