// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2026 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

// Test error when case matches is used with non-tagged union type

module t;
  // Regular union (not tagged)
  union packed {
    int a;
    int b;
  } u;

  initial begin
    // verilator lint_off WIDTHEXPAND
    case (u) matches
      tagged Valid .v: $display("valid");
      default: $display("default");
    endcase
    // verilator lint_on WIDTHEXPAND
  end
endmodule
