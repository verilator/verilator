// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2022 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

extern program ex_pgm;
extern interface ex_ifc;
extern module ex_mod;

module t;

  ex_pgm u_pgm();
  ex_ifc u_ifc();
  ex_mod u_mod();

  initial begin
    $write("*-* All Finished *-*\n");
    $finish;
  end

endmodule

// Could be in another compile run, but we don't support that
program ex_pgm;
endprogram

interface ex_ifc;
endinterface

module ex_mod;
endmodule
