// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2020 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

class Cls;
   function void pre_randomize;
   endfunction;

   function void post_randomize;
   endfunction;
endclass

module t (/*AUTOARG*/);
endmodule
