// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2009 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;
   reg foobar;

   task boobar; endtask

   initial begin
      if (foobat) $stop;
      boobat;
   end
endmodule
