module t;
endmodule
