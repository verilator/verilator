// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2016 by Wilson Snyder.

module t (/*AUTOARG*/);

   shortreal s;

   initial s = 1.2345;

endmodule
