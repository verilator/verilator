// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2023 Antmicro Ltd
// SPDX-License-Identifier: CC0-1.0

class Bar#(type T = int);
   T t;
   function new;
      t = new;
   endfunction
endclass

class Baz;
   int x = 1;
endclass

module t;
   initial begin
      Bar#(Baz) bar_baz = new;
      if (bar_baz.t.x != 1) $stop;

      $write("*-* All Finished *-*\n");
      $finish;
   end
endmodule
