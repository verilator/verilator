// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2019 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

virtual class VBase;
endclass

module t;
   initial begin
      automatic VBase b = new;  // Error
   end
endmodule
