// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2023 Antmicro Ltd
// SPDX-License-Identifier: CC0-1.0

module t;

   class bar #(type T) extends T;
   endclass

   typedef real real_t;

   bar #(real_t) bar_real_t;

   initial begin
      $stop;
   end
endmodule
