// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2023 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;
   sub s1();
endmodule

module sub;
   enum {s0, s1} state;
   initial begin
      $write("*-* All Finished *-*\n");
      $finish;
   end
endmodule
