// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2024 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

virtual class Base;
    pure constraint raint;
endclass

class Cls extends Base;
   // Bad: Missing 'constraint raint'
endclass

module t;
endmodule
