// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2010 by Wilson Snyder.

module t;
   t_lint_declfilename sub ();
endmodule

module t_lint_declfilename;
endmodule
