// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain.
// SPDX-FileCopyrightText: 2025 Wilson Snyder
// SPDX-License-Identifier: CC0-1.0

module t;

  bit bad = '{1'b1};  // <--- BAD: Can't assign pattern to scalar

  initial $stop;
endmodule
