// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2025 by Antmicro.
// SPDX-License-Identifier: CC0-1.0

/* verilator lint_off COVERIGN */
module t();
    covergroup cg;
    function sample();

    endfunction
    function get_coverage();

    endfunction
    endgroup
endmodule
